`define LDM_DEPTH 8
`define CTX_RC_DEPTH 2960
`define CTX_PE_DEPTH 2960
`define CTX_IM_DEPTH 2960
