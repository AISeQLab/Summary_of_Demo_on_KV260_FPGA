`define LDM_DEPTH 32
`define CTX_RC_DEPTH 192
`define CTX_PE_DEPTH 192
`define CTX_IM_DEPTH 192
