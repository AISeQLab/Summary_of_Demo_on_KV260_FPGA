`define LDM_DEPTH 48
`define CTX_RC_DEPTH 1060
`define CTX_PE_DEPTH 1060
`define CTX_IM_DEPTH 1060
