`define LDM_DEPTH 32
`define CTX_RC_DEPTH 432
`define CTX_PE_DEPTH 432
`define CTX_IM_DEPTH 432
