`define LDM_DEPTH 32
`define CTX_RC_DEPTH 11552
`define CTX_PE_DEPTH 11552
`define CTX_IM_DEPTH 11552
