`define LDM_DEPTH 32
`define CTX_RC_DEPTH 672
`define CTX_PE_DEPTH 672
`define CTX_IM_DEPTH 672
